`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:34:38 12/16/2018 
// Design Name: 
// Module Name:    Clock12MergedDispDecoder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Clock12MergedDispDecoder(
	input is_on,
	
	// set related
	input [1:0] current_set_state,
	input set_isPM 
    );


endmodule
